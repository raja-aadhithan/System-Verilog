interface intf();
  logic [3:0] a,b,sum;
  logic cy;
endinterface