interface intf();
  logic a,b,sum,carry;
endinterface